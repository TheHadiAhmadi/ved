module main 

import editor

fn main() {
    editor.initialize()
}
